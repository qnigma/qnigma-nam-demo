localparam REFCLK_HZ = 125000000;